* circuit testbench

* Include the specific transistor models
.lib "/usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* Include the mux2_1 subcircuit
.include mux2_1.mod

ahdldevice [clock reset] [d0 d1 s] null dmod VHI=1.8 VLO=0
.model dmod d_cosim simulation "./stim_gen.so"* Instantiate mux

X0 d0 d1 s y mux2_1

* Clock generator
Vclock clock 0 PULSE(0 1.8 0 1n 1n 10n 20n)
Vreset reset 0 PULSE(0 1.8 0 1n 1n 10n 0)

.control

  tran 1n 200n
  plot v(d0) 
  plot v(d1) 
  plot v(s) 
  plot v(y)

.endc


.end
